module main(); endmodule